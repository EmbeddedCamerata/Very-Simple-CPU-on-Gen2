`define INS_LENGTH 	4

`define REG_NUM		4
`define CODE_WIDTH	2

`define CMD_LENGTH 	6
`define CMD_MV 		(2'b00)
`define CMD_MVI 	(2'b01)
`define CMD_ADD 	(2'b10)
`define CMD_SUB 	(2'b11)

`define ALU_ADD		(1'b0)
`define ALU_SUB		(1'b1)